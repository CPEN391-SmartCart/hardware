module Path_Writer(
	input logic clk,
	input logic reset,


);


	enum logic [2:0] {
		IDLE,
		START,

	} state;

	

endmodule